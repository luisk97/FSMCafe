module Expreso ()