module agua (output logic s);

	assign s = 1;
endmodule;