module agua (input logic i, output logic s);

	assign s = i;
endmodule 