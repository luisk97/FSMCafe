module cafe (output logic s);

	assign s = 1'b1;

endmodule